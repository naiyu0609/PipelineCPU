module Adder(
 	input [31:0] data1,//Number1
 	input [31:0] data2,//Number2
 	output [31:0] data_o//Result
);

assign data_o=data1+data2;//Function

endmodule
